module stopwatch(
    input clk,
    input mod, //если 0 значит режим секундомера
    input key_start,
    input key_reset,

    output logic [3:0] Hex_0,
    output logic [3:0] Hex_1,
    output logic [3:0] Hex_2,
    output logic [3:0] Hex_3
);
localparam  IN_CLK_HZ = 50_000_000;
localparam  MM_count=IN_CLK_HZ/100;

typedef enum logic[1:0] {SHOW_MM, SHOW_SS} show_t;

show_t show_next, show_state;

logic [25:0] count = 1;

logic start_stop ='0;

logic [3:0] time_S  =0;
logic [3:0] time_SS =0;
logic [3:0] time_M  =0;
logic [3:0] time_MM =0;

always_comb begin
	show_next = SHOW_MM;
    case (show_state)
    SHOW_MM:
        if ((time_MM >=5) && (time_M >=4'b1001) && (time_SS >=4'b1001) && (time_S >=4'b1001) && (count >= MM_count))
            show_next = SHOW_SS;
        else
            show_next = SHOW_MM;
    SHOW_SS: show_next = SHOW_SS;
    default: show_next = SHOW_MM;    
    endcase
end

always_ff @(posedge clk or posedge key_reset)
    if (!mod) begin
        if (key_reset)
            show_state <= SHOW_MM;
        else
            show_state <= show_next;
    end

always_ff@(posedge clk) begin
    if(!mod) begin
        Hex_0 <= time_S;
        Hex_1 <= time_SS;
        Hex_2 <= time_M;
        Hex_3 <= time_MM;
    end
end    
//----------------------------------------------------------------------------//
always_ff @(posedge clk or posedge key_reset)
    if(!mod) begin
        if (key_reset) begin
            time_S  <= 0;
            time_SS <= 0;
            time_M  <= 0;
            time_MM <= 0;   
            start_stop <= '0;
        end
        else begin
            if (key_start) 
                start_stop <= ~start_stop;                  
            
            if (start_stop)                
                count <= count +1'b1;

            case (show_state)
            SHOW_MM: SS_MM();
            SHOW_SS: MM_SS();
            default: MM_SS();
            endcase                             
        end
    end
//-------------------------------------------------------------------------//
task SS_MM();
       if (count >= MM_count) begin                        
            if (time_S >=4'b1001) begin               
                time_S  <= 4'b0000;
                if (time_SS >=4'b1001) begin 
                    time_SS <= 4'b0000;
                   if (time_M >=4'b1001) begin 
                       time_M <= 4'b0000;
                       if (time_MM >=5) begin 
                           time_MM <= 4'b0000;
                           time_M  <= 4'b0001;
                           time_SS <= 4'b0000;
                           time_S  <= 4'b0000;
                       end else 
                           time_MM <= time_MM +1'b1;
                    end else 
                        time_M <= time_M +1'b1;
                end else 
                    time_SS <= time_SS+4'b0001;
            end else          
                time_S <= time_S+1'b1;
            count <= '0;
        end         
    endtask : SS_MM
//------------------------------------------------------------------------//
task MM_SS();        
        if (count >= IN_CLK_HZ) begin                        
            if (time_S==4'b1001) begin               
                time_S  <= 4'b0000;
                if (time_SS==4'b0101) begin 
                    time_SS <= 4'b0000;
                   if (time_M==4'b1001) begin 
                       time_M <= 4'b0000;
                       if (time_MM==4'b0101) begin 
                           time_MM <= 4'b0000;
                           time_M  <= 4'b0000;
                           time_SS <= 4'b0000;
                           time_M  <= 4'b0000;
                       end else 
                           time_MM <= time_MM +1'b1;
                    end else 
                        time_M <= time_M +1'b1;
                end else 
                    time_SS <= time_SS+1'b1;
            end else          
                time_S <= time_S+1'b1;
            count <= '0;
        end          
    endtask : MM_SS
    //---------------------------------------------------------------------------//	 
//------------------------------------------------------------------------//
endmodule :stopwatch